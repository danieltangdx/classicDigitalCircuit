/******************
	FileName	:	decodeThreetoEight.v
	Author		:	daniel
	Description	:	Example of a 3-8 decode
	Revision	:	2017/12/20
	Company		:	***********
	code		:	Verilog-2001
************************/
module decodeThreeoEight(
input 					iEnable,
input				[2:0]	iA,
output	reg	[7:0]	oA);
always @(iEnable or iA)
begin
	if(!iEnable)
		oA = 8'b0;
	else
		case(iA)
		3'b000: oA = 8'b0000_0001;
		3'b001: oA = 8'b0000_0010;
		3'b010: oA = 8'b0000_0100;
		3'b011: oA = 8'b0000_1000;
		3'b100: oA = 8'b0001_0000;
		3'b101: oA = 8'b0010_0000;
		3'b110: oA = 8'b0100_0000;
		3'b111: oA = 8'b1000_0000;
		default:oA = 8'b0000_0000;
		endcase
end
endmodule
